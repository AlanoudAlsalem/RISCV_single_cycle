module control_unit #(
    `include "parameters.vh"
)(
    input   [6:0] opcode,
    input   [2:0] funct3,
    input   [6:0] funct7,
);

endmodule