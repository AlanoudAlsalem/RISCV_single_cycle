parameter
// op codes                     // funct3               // funct7
lb_op       =   7'b0000011,     lb_f3   =   3'b000,     
lh_op       =   7'b0000011,     lh_f3   =   3'b001,
lw_op       =   7'b0000011,     lw_f3   =   3'b010,
ld_op       =   7'b0000011,     lf_f3   =   3'b011,
lbu_op      =   7'b0000011,     lbu_f3  =   3'b100,
lhu_op      =   7'b0000011,     lhu_f3  =   3'b101,
lwu_op      =   7'b0000011,     lwu_f3  =   3'b110,
addi_op     =   7'b0010011,     addi_f3 =   3'b000,
slli_op     =   7'b0010011,     slli_f3 =   3'b001,     slli_f7 =   7'b0000000,   
slti_op     =   7'b0010011,     slti_f3 =   3'b010,
xori_op     =   7'b0010011,     xori_f3 =   3'b100,
srli_op     =   7'b0010011,     srli_f3 =   3'b101,     srli_f7 =   7'b0000000,
ori_op      =   7'b0010011,     ori_f3  =   3'b110,
andi_op     =   7'b0010011,     andi_f3 =   3'b111,   
sb_op       =   7'b0100011,     sb_f3   =   3'b000,
sw_op       =   7'b0100011,     sw_f3   =   3'b010,
add_op      =   7'b0110011,     add_f3  =   3'b000,     add_f7  =   7'b0000000,  
sub_op      =   7'b0110011,     sub_f3  =   3'b000,     sub_f7  =   7'b0100000,
sll_op      =   7'b0110011,     sll_f3  =   3'b001,     sll_f7  =   7'b0000000,
slt_op      =   7'b0110011,     slt_f3  =   3'b010,     slt_f7  =   7'b0000000,
xor_op      =   7'b0110011,     xor_f3  =   3'b100,     xor_f6  =   7'b0000000,
srl_op      =   7'b0110011,     srl_f3  =   3'b101,     srl_f7  =   7'b0000000,
or_op       =   7'b0110011,     or_f3   =   3'b110,     or_f7   =   7'b0000000,
and_op      =   7'b0110011,     and_f3  =   3'b111,     and_f7  =   7'b0000000,
lui_op      =   7'b0110111,
beq_op      =   7'b1100011,     beq_f3  =   3'b000,
bne_op      =   7'b1100011,     bne_f3  =   3'b001,
blt_op      =   7'b1100011,     blt_f3  =   3'b100,
bge_op      =   7'b1100011,     bge_f3  =   3'b101,
jalr_op     =   7'b1100111,     jalr_f3 =   3'b000,
jal_op      =   7'b1101111,

//ALU operations
add_    = 4'b0001,
sub_    = 4'b0010,
and_    = 4'b0011,
or_     = 4'b0100,
sll_    = 4'b0101,
srl_    = 4'b0110,
xor_    = 4'b0111,
slt_    = 4'b1000,
jal_    = 4'b1001,
lui_    = 4'b1010